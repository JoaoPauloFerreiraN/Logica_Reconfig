library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all

entity barrelShifter is
	generic (N: integer :=4);
	port (a: in std_logic_vector (N-1 downto 0);
			s: out std_logic_vector (N-1 downto 0));
end entity;

architecture arq of barrelShifter is
	type vec_int is array (N-1 downto 0) of integer range 0 to N;
	signal vecAux, vecAux2: vec_int;
	begin
	
	vecAux(to_integer(unsigned(a))) <= a;	
	gen_1: for i in 0 to N-1 generate
		vecAux2(i) <=( others => '0'); -- cria vetor de zeros
	end generate;
		
		gen_2: for j in 0 to N-1 generate
			if 
	
	
	
	
end architecture;
	